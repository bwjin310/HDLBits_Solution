module top_module (
    input [3:0] SW, //R
    input [3:0] KEY, //w, L, E
    output [3:0] LEDR //output
); //注意接口顺序

    mux2_Dff ins1(
        .clk(KEY[0]),
        .w(KEY[3]),
        .R(SW[3]),
        .E(KEY[1]),
        .L(KEY[2]),
        .Q(LEDR[3])
    );
    mux2_Dff ins2(
        .clk(KEY[0]),
        .w(LEDR[3]),
        .R(SW[2]),
        .E(KEY[1]),
        .L(KEY[2]),
        .Q(LEDR[2])
    );
    mux2_Dff ins3(
        .clk(KEY[0]),
        .w(LEDR[2]),
        .R(SW[1]),
        .E(KEY[1]),
        .L(KEY[2]),
        .Q(LEDR[1])
    );
    mux2_Dff ins4(
        .clk(KEY[0]),
        .w(LEDR[1]),
        .R(SW[0]),
        .E(KEY[1]),
        .L(KEY[2]),
        .Q(LEDR[0])
    );
endmodule

module mux2_Dff (
    input clk,
    input w, R, E, L,
    output Q
);

    always @(posedge clk ) begin
        Q <= L? R : E? w : Q;
    end
endmodule