module top_module (
    input clk,
    input enable,
    input S,
    input A, B, C,
    output Z ); 

endmodule
