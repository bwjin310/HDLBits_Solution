module top_module (
    output zero // no colon after word output
);
    assign zero = 1'b0;
endmodule
